/**
 * @file	InstMem.vh
 * @author	LiuChuanXi
 * @date	2021.04.28
 * @version	V1.0
 * @brief	InstMem模块的宏定义
 * @par	修改日志
 * <table>
 * <tr><th>Date			<th>Version		<th>Author		<th>Description
 * <tr><td>2021.04.28	<td>V1.0		<td>LiuChuanXi	<td>创建初始版本
 * </table>
 */

`ifndef __INSTMEM_H
`define __INSTMEM_H

/* ROM的长和宽，以及地址位数 */
`define WIDTH_ROM		8		//width of the rom
`define DEPTH_ROM		256		//depth of the rom
`define LEN_ADDR_ROM	8		//length of the rom address


`endif // __INSTMEM_H
